library verilog;
use verilog.vl_types.all;
entity Lab04_vlg_vec_tst is
end Lab04_vlg_vec_tst;
