library verilog;
use verilog.vl_types.all;
entity MUX8bit_vlg_vec_tst is
end MUX8bit_vlg_vec_tst;
