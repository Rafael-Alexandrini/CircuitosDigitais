library verilog;
use verilog.vl_types.all;
entity cla_vlg_vec_tst is
end cla_vlg_vec_tst;
